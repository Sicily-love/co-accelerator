module PE_array1#(
    parameter WORDWIDTH = 32
)
(

);


endmodule